--
--
--
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity A429_Tx is
    generic();
    port();
end entity;

architecture main of A429_Tx is
begin
end architecture;